`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Alex Buhse
// 
// Create Date:    21:21:22 12/03/2016 
// Design Name: 
// Module Name:    EksBlowfishSetup 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module EksBlowfishSetup(
    input clk,
    input [127:0] Salt,
    input [7:0] cost,
    input [575:0] Key,
	 input rst,
    output[327:0] cryptm
    );
	 
	 integer j;
	 integer i;
	 integer q;
	 integer y;
	 integer ecb;
	 reg initDone;
	 reg expandDone;
	 reg [191:0] cyph;
	 reg [63:0] ctext;
	 reg [31:0] P [0:17];
	 reg [31:0] S0 [0:255];
	 reg [31:0] S1 [0:255];
	 reg [31:0] S2 [0:255];
	 reg [31:0] S3 [0:255];
	 reg [327:0] cryptmw;
	 
	function [31:0] f;
	input [31:0] inp;
	reg [31:0] t0;
	reg [31:0] t1;
	begin
	f = S0[inp[31:24]] + S1[inp[23:16]];
	f = f ^ S2[inp[15:8]] + S3[inp[7:0]];
	//f = t1 + S3[inp[7:0]];
	end
	endfunction
	
	function [63:0] Encrypt;
	input [63:0] sal;
	reg [31:0] l;
	reg [31:0] r;
	reg [31:0] temp;
	begin
	l = sal[63:32];
	r = sal[31:0];
	for(i = 0; i < 16; i = i + 2)
		begin
		l = l ^ P[i];
		r = r ^ f(l);
		r = r ^ P[i + 1];
		l = l ^ f(r);
		end
	l = l ^ P[16];
	r = r ^ P[17];
	temp = r;
	r = l;
	l = temp;
	Encrypt = {l,r};
	end
	endfunction
	
	task expandKey;
	input [127:0] salt;
	input [575:0] key;
		begin
		P[0] = key[575:544] ^ P[0];
		P[1] = key[543:512] ^ P[1];
		P[2] = key[511:480] ^ P[2];
		P[3] = key[479:448] ^ P[3];
		P[4] = key[447:416] ^ P[4];
		P[5] = key[415:384] ^ P[5];
		P[6] = key[383:352] ^ P[6];
		P[7] = key[351:320] ^ P[7];
		P[8] = key[319:288] ^ P[8];
		P[9] = key[287:256] ^ P[9];
		P[10] = key[255:224] ^ P[10];
		P[11] = key[223:192] ^ P[11];
		P[12] = key[191:160] ^ P[12];
		P[13] = key[159:128] ^ P[13];
		P[14] = key[127:96] ^ P[14];
		P[15] = key[95:64] ^ P[15];
		P[16] = key[63:32] ^ P[16];
		P[17] = key[31:0] ^ P[17];

		ctext = Encrypt(salt[127:64]);

		P[0] = ctext[63:32];
		P[1] = ctext[31:0];

		//n = 2
		ctext = Encrypt(ctext ^ salt[127:64]);
		P[2] = ctext[63:32];
		P[3] = ctext[31:0];
		
		//n = 3
		ctext = Encrypt(ctext ^ salt[63:0]);
		P[4] = ctext[63:32];
		P[5] = ctext[31:0];

		//n = 4
		ctext = Encrypt(ctext ^ salt[127:64]);
		P[6] = ctext[63:32];
		P[7] = ctext[31:0];

		//n = 5
		ctext = Encrypt(ctext ^ salt[63:0]);
		P[8] = ctext[63:32];
		P[9] = ctext[31:0];

		//n = 6
		ctext = Encrypt(ctext ^ salt[127:64]);
		P[10] = ctext[63:32];
		P[11] = ctext[31:0];

		//n = 7
		ctext = Encrypt(ctext ^ salt[63:0]);
		P[12] = ctext[63:32];
		P[13] = ctext[31:0];

		//n = 8
		ctext = Encrypt(ctext ^ salt[127:64]);
		P[14] = ctext[63:32];
		P[15] = ctext[31:0];

		//n = 9
		ctext = Encrypt(ctext ^ salt[63:0]);
		P[16] = ctext[63:32];
		P[17] = ctext[31:0];
		
		for (j = 0; j < 64; j = j + 4)
			begin
			ctext = Encrypt(ctext ^ salt[127:64]);
			S0[4 * j] = ctext[63:32];
			S0[4 * j + 1] = ctext[31:0];
			ctext = Encrypt(ctext ^ salt[63:0]);
			S0[4 * j + 2] = ctext[63:32];
			S0[4 * j + 3] = ctext[31:0];
			end
		
		for (j = 0; j < 64; j = j + 4)
			begin
			ctext = Encrypt(ctext ^ salt[127:64]);
			S1[4 * j] = ctext[63:32];
			S1[4 * j + 1] = ctext[31:0];
			ctext = Encrypt(ctext ^ salt[63:0]);
			S1[4 * j + 2] = ctext[63:32];
			S1[4 * j + 3] = ctext[31:0];
			end
		
		for (j = 0; j < 64; j = j + 4)
			begin
			ctext = Encrypt(ctext ^ salt[127:64]);
			S2[4 * j] = ctext[63:32];
			S2[4 * j + 1] = ctext[31:0];
			ctext = Encrypt(ctext ^ salt[63:0]);
			S2[4 * j + 2] = ctext[63:32];
			S2[4 * j + 3] = ctext[31:0];
			end
		
		for (j = 0; j < 64; j = j + 4)
			begin
			ctext = Encrypt(ctext ^ salt[127:64]);
			S3[4 * j] = ctext[63:32];
			S3[4 * j + 1] = ctext[31:0];
			ctext = Encrypt(ctext ^ salt[63:0]);
			S3[4 * j + 2] = ctext[63:32];
			S3[4 * j + 3] = ctext[31:0];
			end
		end
		
	endtask
	 
	 always @(posedge clk, posedge rst)
	begin
	 
		if(rst)
		begin
			
			initDone = 0;
			expandDone = 0;
			P[0] <= 32'h243f6a88;
			P[1] <= 32'h85a308d3;
			P[2] <= 32'h13198a2e;
			P[3] <= 32'h03707344;
			P[4] <= 32'ha4093822;
			P[5] <= 32'h299f31d0;
			P[6] <= 32'h082efa98;
			P[7] <= 32'hec4e6c89;
			P[8] <= 32'h452821e6;
			P[9] <= 32'h38d01377;
			P[10] <= 32'hbe5466cf;
			P[11] <= 32'h34e90c6c;
			P[12] <= 32'hc0ac29b7;
			P[13] <= 32'hc97c50dd;
			P[14] <= 32'h3f84d5b5;
			P[15] <= 32'hb5470917;
			P[16] <= 32'h9216d5d9;
			P[17] <= 32'h8979fb1b;
			
			cyph <= 192'h4f72706865616e4265686f6c64657253637279446f756274;
			
			
			S0[0] <= 32'hd1310ba6; S0[1] <= 32'h98dfb5ac; S0[2] <= 32'h2ffd72db;
			S0[3] <= 32'hd01adfb7; S0[4] <= 32'hb8e1afed; S0[5] <= 32'h6a267e96;
			S0[6] <= 32'hba7c9045; S0[7] <= 32'hf12c7f99; S0[8] <= 32'h24a19947;
			S0[9] <= 32'hb3916cf7; S0[10] <= 32'h0801f2e2; S0[11] <= 32'h858efc16;
			S0[12] <= 32'h636920d8; S0[13] <= 32'h71574e69; S0[14] <= 32'ha458fea3;
			S0[15] <= 32'hf4933d7e; S0[16] <= 32'h0d95748f; S0[17] <= 32'h728eb658;
			S0[18] <= 32'h718bcd58; S0[19] <= 32'h82154aee; S0[20] <= 32'h7b54a41d;
			S0[21] <= 32'hc25a59b5; S0[22] <= 32'h9c30d539; S0[23] <= 32'h2af26013;
			S0[24] <= 32'hc5d1b023; S0[25] <= 32'h286085f0; S0[26] <= 32'hca417918;
			S0[27] <= 32'hb8db38ef; S0[28] <= 32'h8e79dcb0; S0[29] <= 32'h603a180e;
			S0[30] <= 32'h6c9e0e8b; S0[31] <= 32'hb01e8a3e; S0[32] <= 32'hd71577c1;
			S0[33] <= 32'hbd314b27; S0[34] <= 32'h78af2fda; S0[35] <= 32'h55605c60;
			S0[36] <= 32'he65525f3; S0[37] <= 32'haa55ab94; S0[38] <= 32'h57489862;
			S0[39] <= 32'h63e81440; S0[40] <= 32'h55ca396a; S0[41] <= 32'h2aab10b6;
			S0[42] <= 32'hb4cc5c34; S0[43] <= 32'h1141e8ce; S0[44] <= 32'ha15486af;
			S0[45] <= 32'h7c72e993; S0[46] <= 32'hb3ee1411; S0[47] <= 32'h636fbc2a;
			S0[48] <= 32'h2ba9c55d; S0[49] <= 32'h741831f6; S0[50] <= 32'hce5c3e16;
			S0[51] <= 32'h9b87931e; S0[52] <= 32'hafd6ba33; S0[53] <= 32'h6c24cf5c;
			S0[54] <= 32'h7a325381; S0[55] <= 32'h28958677; S0[56] <= 32'h3b8f4898;
			S0[57] <= 32'h6b4bb9af; S0[58] <= 32'hc4bfe81b; S0[59] <= 32'h66282193;
			S0[60] <= 32'h61d809cc; S0[61] <= 32'hfb21a991; S0[62] <= 32'h487cac60;
			S0[63] <= 32'h5dec8032; S0[64] <= 32'hef845d5d; S0[65] <= 32'he98575b1;
			S0[66] <= 32'hdc262302; S0[67] <= 32'heb651b88; S0[68] <= 32'h23893e81;
			S0[69] <= 32'hd396acc5; S0[70] <= 32'h0f6d6ff3; S0[71] <= 32'h83f44239;
			S0[72] <= 32'h2e0b4482; S0[73] <= 32'ha4842004; S0[74] <= 32'h69c8f04a;
			S0[75] <= 32'h9e1f9b5e; S0[76] <= 32'h21c66842; S0[77] <= 32'hf6e96c9a;
			S0[78] <= 32'h670c9c61; S0[79] <= 32'habd388f0; S0[80] <= 32'h6a51a0d2;
			S0[81] <= 32'hd8542f68; S0[82] <= 32'h960fa728; S0[83] <= 32'hab5133a3;
			S0[84] <= 32'h6eef0b6c; S0[85] <= 32'h137a3be4; S0[86] <= 32'hba3bf050;
			S0[87] <= 32'h7efb2a98; S0[88] <= 32'ha1f1651d; S0[89] <= 32'h39af0176;
			S0[90] <= 32'h66ca593e; S0[91] <= 32'h82430e88; S0[92] <= 32'h8cee8619;
			S0[93] <= 32'h456f9fb4; S0[94] <= 32'h7d84a5c3; S0[95] <= 32'h3b8b5ebe;
			S0[96] <= 32'he06f75d8; S0[97] <= 32'h85c12073; S0[98] <= 32'h401a449f;
			S0[99] <= 32'h56c16aa6; S0[100] <= 32'h4ed3aa62; S0[101] <= 32'h363f7706;
			S0[102] <= 32'h1bfedf72; S0[103] <= 32'h429b023d; S0[104] <= 32'h37d0d724;
			S0[105] <= 32'hd00a1248; S0[106] <= 32'hdb0fead3; S0[107] <= 32'h49f1c09b;
			S0[108] <= 32'h075372c9; S0[109] <= 32'h80991b7b; S0[110] <= 32'h25d479d8;
			S0[111] <= 32'hf6e8def7; S0[112] <= 32'he3fe501a; S0[113] <= 32'hb6794c3b;
			S0[114] <= 32'h976ce0bd; S0[115] <= 32'h04c006ba; S0[116] <= 32'hc1a94fb6;
			S0[117] <= 32'h409f60c4; S0[118] <= 32'h5e5c9ec2; S0[119] <= 32'h196a2463;
			S0[120] <= 32'h68fb6faf; S0[121] <= 32'h3e6c53b5; S0[122] <= 32'h1339b2eb;
			S0[123] <= 32'h3b52ec6f; S0[124] <= 32'h6dfc511f; S0[125] <= 32'h9b30952c;
			S0[126] <= 32'hcc814544; S0[127] <= 32'haf5ebd09; S0[128] <= 32'hbee3d004;
			S0[129] <= 32'hde334afd; S0[130] <= 32'h660f2807; S0[131] <= 32'h192e4bb3;
			S0[132] <= 32'hc0cba857; S0[133] <= 32'h45c8740f; S0[134] <= 32'hd20b5f39;
			S0[135] <= 32'hb9d3fbdb; S0[136] <= 32'h5579c0bd; S0[137] <= 32'h1a60320a;
			S0[138] <= 32'hd6a100c6; S0[139] <= 32'h402c7279; S0[140] <= 32'h679f25fe;
			S0[141] <= 32'hfb1fa3cc; S0[142] <= 32'h8ea5e9f8; S0[143] <= 32'hdb3222f8;
			S0[144] <= 32'h3c7516df; S0[145] <= 32'hfd616b15; S0[146] <= 32'h2f501ec8;
			S0[147] <= 32'had0552ab; S0[148] <= 32'h323db5fa; S0[149] <= 32'hfd238760;
			S0[150] <= 32'h53317b48; S0[151] <= 32'h3e00df82; S0[152] <= 32'h9e5c57bb;
			S0[153] <= 32'hca6f8ca0; S0[154] <= 32'h1a87562e; S0[155] <= 32'hdf1769db;
			S0[156] <= 32'hd542a8f6; S0[157] <= 32'h287effc3; S0[158] <= 32'hac6732c6;
			S0[159] <= 32'h8c4f5573; S0[160] <= 32'h695b27b0; S0[161] <= 32'hbbca58c8;
			S0[162] <= 32'he1ffa35d; S0[163] <= 32'hb8f011a0; S0[164] <= 32'h10fa3d98;
			S0[165] <= 32'hfd2183b8; S0[166] <= 32'h4afcb56c; S0[167] <= 32'h2dd1d35b;
			S0[168] <= 32'h9a53e479; S0[169] <= 32'hb6f84565; S0[170] <= 32'hd28e49bc;
			S0[171] <= 32'h4bfb9790; S0[172] <= 32'he1ddf2da; S0[173] <= 32'ha4cb7e33;
			S0[174] <= 32'h62fb1341; S0[175] <= 32'hcee4c6e8; S0[176] <= 32'hef20cada;
			S0[177] <= 32'h36774c01; S0[178] <= 32'hd07e9efe; S0[179] <= 32'h2bf11fb4;
			S0[180] <= 32'h95dbda4d; S0[181] <= 32'hae909198; S0[182] <= 32'heaad8e71;
			S0[183] <= 32'h6b93d5a0; S0[184] <= 32'hd08ed1d0; S0[185] <= 32'hafc725e0;
			S0[186] <= 32'h8e3c5b2f; S0[187] <= 32'h8e7594b7; S0[188] <= 32'h8ff6e2fb;
			S0[189] <= 32'hf2122b64; S0[190] <= 32'h8888b812; S0[191] <= 32'h900df01c;
			S0[192] <= 32'h4fad5ea0; S0[193] <= 32'h688fc31c; S0[194] <= 32'hd1cff191;
			S0[195] <= 32'hb3a8c1ad; S0[196] <= 32'h2f2f2218; S0[197] <= 32'hbe0e1777;
			S0[198] <= 32'hea752dfe; S0[199] <= 32'h8b021fa1; S0[200] <= 32'he5a0cc0f;
			S0[201] <= 32'hb56f74e8; S0[202] <= 32'h18acf3d6; S0[203] <= 32'hce89e299;
			S0[204] <= 32'hb4a84fe0; S0[205] <= 32'hfd13e0b7; S0[206] <= 32'h7cc43b81;
			S0[207] <= 32'hd2ada8d9; S0[208] <= 32'h165fa266; S0[209] <= 32'h80957705;
			S0[210] <= 32'h93cc7314; S0[211] <= 32'h211a1477; S0[212] <= 32'he6ad2065;
			S0[213] <= 32'h77b5fa86; S0[214] <= 32'hc75442f5; S0[215] <= 32'hfb9d35cf;
			S0[216] <= 32'hebcdaf0c; S0[217] <= 32'h7b3e89a0; S0[218] <= 32'hd6411bd3;
			S0[219] <= 32'hae1e7e49; S0[220] <= 32'h00250e2d; S0[221] <= 32'h2071b35e;
			S0[222] <= 32'h226800bb; S0[223] <= 32'h57b8e0af; S0[224] <= 32'h2464369b;
			S0[225] <= 32'hf009b91e; S0[226] <= 32'h5563911d; S0[227] <= 32'h59dfa6aa;
			S0[228] <= 32'h78c14389; S0[229] <= 32'hd95a537f; S0[230] <= 32'h207d5ba2;
			S0[231] <= 32'h02e5b9c5; S0[232] <= 32'h83260376; S0[233] <= 32'h6295cfa9;
			S0[234] <= 32'h11c81968; S0[235] <= 32'h4e734a41; S0[236] <= 32'hb3472dca;
			S0[237] <= 32'h7b14a94a; S0[238] <= 32'h1b510052; S0[239] <= 32'h9a532915;
			S0[240] <= 32'hd60f573f; S0[241] <= 32'hbc9bc6e4; S0[242] <= 32'h2b60a476;
			S0[243] <= 32'h81e67400; S0[244] <= 32'h08ba6fb5; S0[245] <= 32'h571be91f;
			S0[246] <= 32'hf296ec6b; S0[247] <= 32'h2a0dd915; S0[248] <= 32'hb6636521;
			S0[249] <= 32'he7b9f9b6; S0[250] <= 32'hff34052e; S0[251] <= 32'hc5855664;
			S0[252] <= 32'h53b02d5d; S0[253] <= 32'ha99f8fa1; S0[254] <= 32'h08ba4799;
			S0[255] <= 32'h6e85076a;
			
			
			S1[0] <= 32'h4b7a70e9; S1[1] <= 32'hb5b32944; S1[2] <= 32'hdb75092e;
			S1[3] <= 32'hc4192623; S1[4] <= 32'had6ea6b0; S1[5] <= 32'h49a7df7d;
			S1[6] <= 32'h9cee60b8; S1[7] <= 32'h8fedb266; S1[8] <= 32'hecaa8c71;
			S1[9] <= 32'h699a17ff; S1[10] <= 32'h5664526c; S1[11] <= 32'hc2b19ee1;
			S1[12] <= 32'h193602a5; S1[13] <= 32'h75094c29; S1[14] <= 32'ha0591340;
			S1[15] <= 32'he4183a3e; S1[16] <= 32'h3f54989a; S1[17] <= 32'h5b429d65;
			S1[18] <= 32'h6b8fe4d6; S1[19] <= 32'h99f73fd6; S1[20] <= 32'ha1d29c07;
			S1[21] <= 32'hefe830f5; S1[22] <= 32'h4d2d38e6; S1[23] <= 32'hf0255dc1;
			S1[24] <= 32'h4cdd2086; S1[25] <= 32'h8470eb26; S1[26] <= 32'h6382e9c6;
			S1[27] <= 32'h021ecc5e; S1[28] <= 32'h09686b3f; S1[29] <= 32'h3ebaefc9;
			S1[30] <= 32'h3c971814; S1[31] <= 32'h6b6a70a1; S1[32] <= 32'h687f3584;
			S1[33] <= 32'h52a0e286; S1[34] <= 32'hb79c5305; S1[35] <= 32'haa500737;
			S1[36] <= 32'h3e07841c; S1[37] <= 32'h7fdeae5c; S1[38] <= 32'h8e7d44ec;
			S1[39] <= 32'h5716f2b8; S1[40] <= 32'hb03ada37; S1[41] <= 32'hf0500c0d;
			S1[42] <= 32'hf01c1f04; S1[43] <= 32'h0200b3ff; S1[44] <= 32'hae0cf51a;
			S1[45] <= 32'h3cb574b2; S1[46] <= 32'h25837a58; S1[47] <= 32'hdc0921bd;
			S1[48] <= 32'hd19113f9; S1[49] <= 32'h7ca92ff6; S1[50] <= 32'h94324773;
			S1[51] <= 32'h22f54701; S1[52] <= 32'h3ae5e581; S1[53] <= 32'h37c2dadc;
			S1[54] <= 32'hc8b57634; S1[55] <= 32'h9af3dda7; S1[56] <= 32'ha9446146;
			S1[57] <= 32'h0fd0030e; S1[58] <= 32'hecc8c73e; S1[59] <= 32'ha4751e41;
			S1[60] <= 32'he238cd99; S1[61] <= 32'h3bea0e2f; S1[62] <= 32'h3280bba1; 
			S1[63] <= 32'h183eb331; S1[64] <= 32'h4e548b38; S1[65] <= 32'h4f6db908;
			S1[66] <= 32'h6f420d03; S1[67] <= 32'hf60a04bf; S1[68] <= 32'h2cb81290; 
			S1[69] <= 32'h24977c79; S1[70] <= 32'h5679b072; S1[71] <= 32'hbcaf89af;
			S1[72] <= 32'hde9a771f; S1[73] <= 32'hd9930810; S1[74] <= 32'hb38bae12; 
			S1[75] <= 32'hdccf3f2e; S1[76] <= 32'h5512721f; S1[77] <= 32'h2e6b7124;
			S1[78] <= 32'h501adde6; S1[79] <= 32'h9f84cd87; S1[80] <= 32'h7a584718; 
			S1[81] <= 32'h7408da17; S1[82] <= 32'hbc9f9abc; S1[83] <= 32'he94b7d8c;
			S1[84] <= 32'hec7aec3a; S1[85] <= 32'hdb851dfa; S1[86] <= 32'h63094366; 
			S1[87] <= 32'hc464c3d2; S1[88] <= 32'hef1c1847; S1[89] <= 32'h3215d908;
			S1[90] <= 32'hdd433b37; S1[91] <= 32'h24c2ba16; S1[92] <= 32'h12a14d43; 
			S1[93] <= 32'h2a65c451; S1[94] <= 32'h50940002; S1[95] <= 32'h133ae4dd;
			S1[96] <= 32'h71dff89e; S1[97] <= 32'h10314e55; S1[98] <= 32'h81ac77d6; 
			S1[99] <= 32'h5f11199b; S1[100] <= 32'h043556f1; S1[101] <= 32'hd7a3c76b;
			S1[102] <= 32'h3c11183b; S1[103] <= 32'h5924a509; S1[104] <= 32'hf28fe6ed; 
			S1[105] <= 32'h97f1fbfa; S1[106] <= 32'h9ebabf2c; S1[107] <= 32'h1e153c6e;
			S1[108] <= 32'h86e34570; S1[109] <= 32'heae96fb1; S1[110] <= 32'h860e5e0a; 
			S1[111] <= 32'h5a3e2ab3; S1[112] <= 32'h771fe71c; S1[113] <= 32'h4e3d06fa;
			S1[114] <= 32'h2965dcb9; S1[115] <= 32'h99e71d0f; S1[116] <= 32'h803e89d6; 
			S1[117] <= 32'h5266c825; S1[118] <= 32'h2e4cc978; S1[119] <= 32'h9c10b36a;
			S1[120] <= 32'hc6150eba; S1[121] <= 32'h94e2ea78; S1[122] <= 32'ha5fc3c53; 
			S1[123] <= 32'h1e0a2df4; S1[124] <= 32'hf2f74ea7; S1[125] <= 32'h361d2b3d;
			S1[126] <= 32'h1939260f; S1[127] <= 32'h19c27960; S1[128] <= 32'h5223a708; 
			S1[129] <= 32'hf71312b6; S1[130] <= 32'hebadfe6e; S1[131] <= 32'heac31f66;
			S1[132] <= 32'he3bc4595; S1[133] <= 32'ha67bc883; S1[134] <= 32'hb17f37d1; 
			S1[135] <= 32'h018cff28; S1[136] <= 32'hc332ddef; S1[137] <= 32'hbe6c5aa5;
			S1[138] <= 32'h65582185; S1[139] <= 32'h68ab9802; S1[140] <= 32'heecea50f; 
			S1[141] <= 32'hdb2f953b; S1[142] <= 32'h2aef7dad; S1[143] <= 32'h5b6e2f84;
			S1[144] <= 32'h1521b628; S1[145] <= 32'h29076170; S1[146] <= 32'hecdd4775; 
			S1[147] <= 32'h619f1510; S1[148] <= 32'h13cca830; S1[149] <= 32'heb61bd96;
			S1[150] <= 32'h0334fe1e; S1[151] <= 32'haa0363cf; S1[152] <= 32'hb5735c90; 
			S1[153] <= 32'h4c70a239; S1[154] <= 32'hd59e9e0b; S1[155] <= 32'hcbaade14;
			S1[156] <= 32'heecc86bc; S1[157] <= 32'h60622ca7; S1[158] <= 32'h9cab5cab; 
			S1[159] <= 32'hb2f3846e; S1[160] <= 32'h648b1eaf; S1[161] <= 32'h19bdf0ca;
			S1[162] <= 32'ha02369b9; S1[163] <= 32'h655abb50; S1[164] <= 32'h40685a32; 
			S1[165] <= 32'h3c2ab4b3; S1[166] <= 32'h319ee9d5; S1[167] <= 32'hc021b8f7;
			S1[168] <= 32'h9b540b19; S1[169] <= 32'h875fa099; S1[170] <= 32'h95f7997e; 
			S1[171] <= 32'h623d7da8; S1[172] <= 32'hf837889a; S1[173] <= 32'h97e32d77;
			S1[174] <= 32'h11ed935f; S1[175] <= 32'h16681281; S1[176] <= 32'h0e358829; 
			S1[177] <= 32'hc7e61fd6; S1[178] <= 32'h96dedfa1; S1[179] <= 32'h7858ba99;
			S1[180] <= 32'h57f584a5; S1[181] <= 32'h1b227263; S1[182] <= 32'h9b83c3ff; 
			S1[183] <= 32'h1ac24696; S1[184] <= 32'hcdb30aeb; S1[185] <= 32'h532e3054;
			S1[186] <= 32'h8fd948e4; S1[187] <= 32'h6dbc3128; S1[188] <= 32'h58ebf2ef; 
			S1[189] <= 32'h34c6ffea; S1[190] <= 32'hfe28ed61; S1[191] <= 32'hee7c3c73;
			S1[192] <= 32'h5d4a14d9; S1[193] <= 32'he864b7e3; S1[194] <= 32'h42105d14; 
			S1[195] <= 32'h203e13e0; S1[196] <= 32'h45eee2b6; S1[197] <= 32'ha3aaabea;
			S1[198] <= 32'hdb6c4f15; S1[199] <= 32'hfacb4fd0; S1[200] <= 32'hc742f442; 
			S1[201] <= 32'hef6abbb5; S1[202] <= 32'h654f3b1d; S1[203] <= 32'h41cd2105;
			S1[204] <= 32'hd81e799e; S1[205] <= 32'h86854dc7; S1[206] <= 32'he44b476a; 
			S1[207] <= 32'h3d816250; S1[208] <= 32'hcf62a1f2; S1[209] <= 32'h5b8d2646;
			S1[210] <= 32'hfc8883a0; S1[211] <= 32'hc1c7b6a3; S1[212] <= 32'h7f1524c3; 
			S1[213] <= 32'h69cb7492; S1[214] <= 32'h47848a0b; S1[215] <= 32'h5692b285;
			S1[216] <= 32'h095bbf00; S1[217] <= 32'had19489d; S1[218] <= 32'h1462b174; 
			S1[219] <= 32'h23820e00; S1[220] <= 32'h58428d2a; S1[221] <= 32'h0c55f5ea;
			S1[222] <= 32'h1dadf43e; S1[223] <= 32'h233f7061; S1[224] <= 32'h3372f092; 
			S1[225] <= 32'h8d937e41; S1[226] <= 32'hd65fecf1; S1[227] <= 32'h6c223bdb;
			S1[228] <= 32'h7cde3759; S1[229] <= 32'hcbee7460; S1[230] <= 32'h4085f2a7; 
			S1[231] <= 32'hce77326e; S1[232] <= 32'ha6078084; S1[233] <= 32'h19f8509e;
			S1[234] <= 32'he8efd855; S1[235] <= 32'h61d99735; S1[236] <= 32'ha969a7aa; 
			S1[237] <= 32'hc50c06c2; S1[238] <= 32'h5a04abfc; S1[239] <= 32'h800bcadc;
			S1[240] <= 32'h9e447a2e; S1[241] <= 32'hc3453484; S1[242] <= 32'hfdd56705;
			S1[243] <= 32'h0e1e9ec9; S1[244] <= 32'hdb73dbd3; S1[245] <= 32'h105588cd;
			S1[246] <= 32'h675fda79; S1[247] <= 32'he3674340; S1[248] <= 32'hc5c43465; 
			S1[249] <= 32'h713e38d8; S1[250] <= 32'h3d28f89e; S1[251] <= 32'hf16dff20;
			S1[252] <= 32'h153e21e7; S1[253] <= 32'h8fb03d4a; S1[254] <= 32'he6e39f2b; 
			S1[255] <= 32'hdb83adf7;


			S2[0] <= 32'he93d5a68; S2[1] <= 32'h948140f7; S2[2] <= 32'hf64c261c; 
			S2[3] <= 32'h94692934; S2[4] <= 32'h411520f7; S2[5] <= 32'h7602d4f7;
			S2[6] <= 32'hbcf46b2e; S2[7] <= 32'hd4a20068; S2[8] <= 32'hd4082471; 
			S2[9] <= 32'h3320f46a; S2[10] <= 32'h43b7d4b7; S2[11] <= 32'h500061af;
			S2[12] <= 32'h1e39f62e; S2[13] <= 32'h97244546; S2[14] <= 32'h14214f74; 
			S2[15] <= 32'hbf8b8840; S2[16] <= 32'h4d95fc1d; S2[17] <= 32'h96b591af;
			S2[18] <= 32'h70f4ddd3; S2[19] <= 32'h66a02f45; S2[20] <= 32'hbfbc09ec; 
			S2[21] <= 32'h03bd9785; S2[22] <= 32'h7fac6dd0; S2[23] <= 32'h31cb8504;
			S2[24] <= 32'h96eb27b3; S2[25] <= 32'h55fd3941; S2[26] <= 32'hda2547e6; 
			S2[27] <= 32'habca0a9a; S2[28] <= 32'h28507825; S2[29] <= 32'h530429f4;
			S2[30] <= 32'h0a2c86da; S2[31] <= 32'he9b66dfb; S2[32] <= 32'h68dc1462; 
			S2[33] <= 32'hd7486900; S2[34] <= 32'h680ec0a4; S2[35] <= 32'h27a18dee;
			S2[36] <= 32'h4f3ffea2; S2[37] <= 32'he887ad8c; S2[38] <= 32'hb58ce006; 
			S2[39] <= 32'h7af4d6b6; S2[40] <= 32'haace1e7c; S2[41] <= 32'hd3375fec;
			S2[42] <= 32'hce78a399; S2[43] <= 32'h406b2a42; S2[44] <= 32'h20fe9e35; 
			S2[45] <= 32'hd9f385b9; S2[46] <= 32'hee39d7ab; S2[47] <= 32'h3b124e8b;
			S2[48] <= 32'h1dc9faf7; S2[49] <= 32'h4b6d1856; S2[50] <= 32'h26a36631; 
			S2[51] <= 32'heae397b2; S2[52] <= 32'h3a6efa74; S2[53] <= 32'hdd5b4332;
			S2[54] <= 32'h6841e7f7; S2[55] <= 32'hca7820fb; S2[56] <= 32'hfb0af54e; 
			S2[57] <= 32'hd8feb397; S2[58] <= 32'h454056ac; S2[59] <= 32'hba489527;
			S2[60] <= 32'h55533a3a; S2[61] <= 32'h20838d87; S2[62] <= 32'hfe6ba9b7; 
			S2[63] <= 32'hd096954b; S2[64] <= 32'h55a867bc; S2[65] <= 32'ha1159a58;
			S2[66] <= 32'hcca92963; S2[67] <= 32'h99e1db33; S2[68] <= 32'ha62a4a56; 
			S2[69] <= 32'h3f3125f9; S2[70] <= 32'h5ef47e1c; S2[71] <= 32'h9029317c;
			S2[72] <= 32'hfdf8e802; S2[73] <= 32'h04272f70; S2[74] <= 32'h80bb155c; 
			S2[75] <= 32'h05282ce3; S2[76] <= 32'h95c11548; S2[77] <= 32'he4c66d22;
			S2[78] <= 32'h48c1133f; S2[79] <= 32'hc70f86dc; S2[80] <= 32'h07f9c9ee; 
			S2[81] <= 32'h41041f0f; S2[82] <= 32'h404779a4; S2[83] <= 32'h5d886e17;
			S2[84] <= 32'h325f51eb; S2[85] <= 32'hd59bc0d1; S2[86] <= 32'hf2bcc18f; 
			S2[87] <= 32'h41113564; S2[88] <= 32'h257b7834; S2[89] <= 32'h602a9c60;
			S2[90] <= 32'hdff8e8a3; S2[91] <= 32'h1f636c1b; S2[92] <= 32'h0e12b4c2; 
			S2[93] <= 32'h02e1329e; S2[94] <= 32'haf664fd1; S2[95] <= 32'hcad18115;
			S2[96] <= 32'h6b2395e0; S2[97] <= 32'h333e92e1; S2[98] <= 32'h3b240b62; 
			S2[99] <= 32'heebeb922; S2[100] <= 32'h85b2a20e; S2[101] <= 32'he6ba0d99;
			S2[102] <= 32'hde720c8c; S2[103] <= 32'h2da2f728; S2[104] <= 32'hd0127845; 
			S2[105] <= 32'h95b794fd; S2[106] <= 32'h647d0862; S2[107] <= 32'he7ccf5f0;
			S2[108] <= 32'h5449a36f; S2[109] <= 32'h877d48fa; S2[110] <= 32'hc39dfd27; 
			S2[111] <= 32'hf33e8d1e; S2[112] <= 32'h0a476341; S2[113] <= 32'h992eff74;
			S2[114] <= 32'h3a6f6eab; S2[115] <= 32'hf4f8fd37; S2[116] <= 32'ha812dc60; 
			S2[117] <= 32'ha1ebddf8; S2[118] <= 32'h991be14c; S2[119] <= 32'hdb6e6b0d;
			S2[120] <= 32'hc67b5510; S2[121] <= 32'h6d672c37; S2[122] <= 32'h2765d43b; 
			S2[123] <= 32'hdcd0e804; S2[124] <= 32'hf1290dc7; S2[125] <= 32'hcc00ffa3;
			S2[126] <= 32'hb5390f92; S2[127] <= 32'h690fed0b; S2[128] <= 32'h667b9ffb; 
			S2[129] <= 32'hcedb7d9c; S2[130] <= 32'ha091cf0b; S2[131] <= 32'hd9155ea3;
			S2[132] <= 32'hbb132f88; S2[133] <= 32'h515bad24; S2[134] <= 32'h7b9479bf; 
			S2[135] <= 32'h763bd6eb; S2[136] <= 32'h37392eb3; S2[137] <= 32'hcc115979;
			S2[138] <= 32'h8026e297; S2[139] <= 32'hf42e312d; S2[140] <= 32'h6842ada7; 
			S2[141] <= 32'hc66a2b3b; S2[142] <= 32'h12754ccc; S2[143] <= 32'h782ef11c;
			S2[144] <= 32'h6a124237; S2[145] <= 32'hb79251e7; S2[146] <= 32'h06a1bbe6; 
			S2[147] <= 32'h4bfb6350; S2[148] <= 32'h1a6b1018; S2[149] <= 32'h11caedfa;
			S2[150] <= 32'h3d25bdd8; S2[151] <= 32'he2e1c3c9; S2[152] <= 32'h44421659; 
			S2[153] <= 32'h0a121386; S2[154] <= 32'hd90cec6e; S2[155] <= 32'hd5abea2a;
			S2[156] <= 32'h64af674e; S2[157] <= 32'hda86a85f; S2[158] <= 32'hbebfe988; 
			S2[159] <= 32'h64e4c3fe; S2[160] <= 32'h9dbc8057; S2[161] <= 32'hf0f7c086;
			S2[162] <= 32'h60787bf8; S2[163] <= 32'h6003604d; S2[164] <= 32'hd1fd8346; 
			S2[165] <= 32'hf6381fb0; S2[166] <= 32'h7745ae04; S2[167] <= 32'hd736fccc;
			S2[168] <= 32'h83426b33; S2[169] <= 32'hf01eab71; S2[170] <= 32'hb0804187; 
			S2[171] <= 32'h3c005e5f; S2[172] <= 32'h77a057be; S2[173] <= 32'hbde8ae24;
			S2[174] <= 32'h55464299; S2[175] <= 32'hbf582e61; S2[176] <= 32'h4e58f48f; 
			S2[177] <= 32'hf2ddfda2; S2[178] <= 32'hf474ef38; S2[179] <= 32'h8789bdc2;
			S2[180] <= 32'h5366f9c3; S2[181] <= 32'hc8b38e74; S2[182] <= 32'hb475f255; 
			S2[183] <= 32'h46fcd9b9; S2[184] <= 32'h7aeb2661; S2[185] <= 32'h8b1ddf84;
			S2[186] <= 32'h846a0e79; S2[187] <= 32'h915f95e2; S2[188] <= 32'h466e598e; 
			S2[189] <= 32'h20b45770; S2[190] <= 32'h8cd55591; S2[191] <= 32'hc902de4c;
			S2[192] <= 32'hb90bace1; S2[193] <= 32'hbb8205d0; S2[194] <= 32'h11a86248; 
			S2[195] <= 32'h7574a99e; S2[196] <= 32'hb77f19b6; S2[197] <= 32'he0a9dc09;
			S2[198] <= 32'h662d09a1; S2[199] <= 32'hc4324633; S2[200] <= 32'he85a1f02; 
			S2[201] <= 32'h09f0be8c; S2[202] <= 32'h4a99a025; S2[203] <= 32'h1d6efe10;
			S2[204] <= 32'h1ab93d1d; S2[205] <= 32'h0ba5a4df; S2[206] <= 32'ha186f20f; 
			S2[207] <= 32'h2868f169; S2[208] <= 32'hdcb7da83; S2[209] <= 32'h573906fe;
			S2[210] <= 32'ha1e2ce9b; S2[211] <= 32'h4fcd7f52; S2[212] <= 32'h50115e01; 
			S2[213] <= 32'ha70683fa; S2[214] <= 32'ha002b5c4; S2[215] <= 32'h0de6d027;
			S2[216] <= 32'h9af88c27; S2[217] <= 32'h773f8641; S2[218] <= 32'hc3604c06; 
			S2[219] <= 32'h61a806b5; S2[220] <= 32'hf0177a28; S2[221] <= 32'hc0f586e0;
			S2[222] <= 32'h006058aa; S2[223] <= 32'h30dc7d62; S2[224] <= 32'h11e69ed7; 
			S2[225] <= 32'h2338ea63; S2[226] <= 32'h53c2dd94; S2[227] <= 32'hc2c21634;
			S2[228] <= 32'hbbcbee56; S2[229] <= 32'h90bcb6de; S2[230] <= 32'hebfc7da1; 
			S2[231] <= 32'hce591d76; S2[232] <= 32'h6f05e409; S2[233] <= 32'h4b7c0188;
			S2[234] <= 32'h39720a3d; S2[235] <= 32'h7c927c24; S2[236] <= 32'h86e3725f; 
			S2[237] <= 32'h724d9db9; S2[238] <= 32'h1ac15bb4; S2[239] <= 32'hd39eb8fc;
			S2[240] <= 32'hed545578; S2[241] <= 32'h08fca5b5; S2[242] <= 32'hd83d7cd3; 
			S2[243] <= 32'h4dad0fc4; S2[244] <= 32'h1e50ef5e; S2[245] <= 32'hb161e6f8;
			S2[246] <= 32'ha28514d9; S2[247] <= 32'h6c51133c; S2[248] <= 32'h6fd5c7e7; 
			S2[249] <= 32'h56e14ec4; S2[250] <= 32'h362abfce; S2[251] <= 32'hddc6c837;
			S2[252] <= 32'hd79a3234; S2[253] <= 32'h92638212; S2[254] <= 32'h670efa8e; 
			S2[255] <= 32'h406000e0;
			
			
			S3[0] <= 32'h3a39ce37; S3[1] <= 32'hd3faf5cf; S3[2] <= 32'habc27737; 
			S3[3] <= 32'h5ac52d1b; S3[4] <= 32'h5cb0679e; S3[5] <= 32'h4fa33742;
			S3[6] <= 32'hd3822740; S3[7] <= 32'h99bc9bbe; S3[8] <= 32'hd5118e9d; 
			S3[9] <= 32'hbf0f7315; S3[10] <= 32'hd62d1c7e; S3[11] <= 32'hc700c47b;
			S3[12] <= 32'hb78c1b6b; S3[13] <= 32'h21a19045; S3[14] <= 32'hb26eb1be; 
			S3[15] <= 32'h6a366eb4; S3[16] <= 32'h5748ab2f; S3[17] <= 32'hbc946e79;
			S3[18] <= 32'hc6a376d2; S3[19] <= 32'h6549c2c8; S3[20] <= 32'h530ff8ee; 
			S3[21] <= 32'h468dde7d; S3[22] <= 32'hd5730a1d; S3[23] <= 32'h4cd04dc6;
			S3[24] <= 32'h2939bbdb; S3[25] <= 32'ha9ba4650; S3[26] <= 32'hac9526e8; 
			S3[27] <= 32'hbe5ee304; S3[28] <= 32'ha1fad5f0; S3[29] <= 32'h6a2d519a;
			S3[30] <= 32'h63ef8ce2; S3[31] <= 32'h9a86ee22; S3[32] <= 32'hc089c2b8; 
			S3[33] <= 32'h43242ef6; S3[34] <= 32'ha51e03aa; S3[35] <= 32'h9cf2d0a4;
			S3[36] <= 32'h83c061ba; S3[37] <= 32'h9be96a4d; S3[38] <= 32'h8fe51550; 
			S3[39] <= 32'hba645bd6; S3[40] <= 32'h2826a2f9; S3[41] <= 32'ha73a3ae1;
			S3[42] <= 32'h4ba99586; S3[43] <= 32'hef5562e9; S3[44] <= 32'hc72fefd3; 
			S3[45] <= 32'hf752f7da; S3[46] <= 32'h3f046f69; S3[47] <= 32'h77fa0a59;
			S3[48] <= 32'h80e4a915; S3[49] <= 32'h87b08601; S3[50] <= 32'h9b09e6ad; 
			S3[51] <= 32'h3b3ee593; S3[52] <= 32'he990fd5a; S3[53] <= 32'h9e34d797;
			S3[54] <= 32'h2cf0b7d9; S3[55] <= 32'h022b8b51; S3[56] <= 32'h96d5ac3a; 
			S3[57] <= 32'h017da67d; S3[58] <= 32'hd1cf3ed6; S3[59] <= 32'h7c7d2d28;
			S3[60] <= 32'h1f9f25cf; S3[61] <= 32'hadf2b89b; S3[62] <= 32'h5ad6b472; 
			S3[63] <= 32'h5a88f54c; S3[64] <= 32'he029ac71; S3[65] <= 32'he019a5e6;
			S3[66] <= 32'h47b0acfd; S3[67] <= 32'hed93fa9b; S3[68] <= 32'he8d3c48d; 
			S3[69] <= 32'h283b57cc; S3[70] <= 32'hf8d56629; S3[71] <= 32'h79132e28;
			S3[72] <= 32'h785f0191; S3[73] <= 32'hed756055; S3[74] <= 32'hf7960e44; 
			S3[75] <= 32'he3d35e8c; S3[76] <= 32'h15056dd4; S3[77] <= 32'h88f46dba;
			S3[78] <= 32'h03a16125; S3[79] <= 32'h0564f0bd; S3[80] <= 32'hc3eb9e15; 
			S3[81] <= 32'h3c9057a2; S3[82] <= 32'h97271aec; S3[83] <= 32'ha93a072a;
			S3[84] <= 32'h1b3f6d9b; S3[85] <= 32'h1e6321f5; S3[86] <= 32'hf59c66fb; 
			S3[87] <= 32'h26dcf319; S3[88] <= 32'h7533d928; S3[89] <= 32'hb155fdf5;
			S3[90] <= 32'h03563482; S3[91] <= 32'h8aba3cbb; S3[92] <= 32'h28517711; 
			S3[93] <= 32'hc20ad9f8; S3[94] <= 32'habcc5167; S3[95] <= 32'hccad925f;
			S3[96] <= 32'h4de81751; S3[97] <= 32'h3830dc8e; S3[98] <= 32'h379d5862; 
			S3[99] <= 32'h9320f991; S3[100] <= 32'hea7a90c2; S3[101] <= 32'hfb3e7bce;
			S3[102] <= 32'h5121ce64; S3[103] <= 32'h774fbe32; S3[104] <= 32'ha8b6e37e; 
			S3[105] <= 32'hc3293d46; S3[106] <= 32'h48de5369; S3[107] <= 32'h6413e680;
			S3[108] <= 32'ha2ae0810; S3[109] <= 32'hdd6db224; S3[110] <= 32'h69852dfd; 
			S3[111] <= 32'h09072166; S3[112] <= 32'hb39a460a; S3[113] <= 32'h6445c0dd;
			S3[114] <= 32'h586cdecf; S3[115] <= 32'h1c20c8ae; S3[116] <= 32'h5bbef7dd; 
			S3[117] <= 32'h1b588d40; S3[118] <= 32'hccd2017f; S3[119] <= 32'h6bb4e3bb;
			S3[120] <= 32'hdda26a7e; S3[121] <= 32'h3a59ff45; S3[122] <= 32'h3e350a44; 
			S3[123] <= 32'hbcb4cdd5; S3[124] <= 32'h72eacea8; S3[125] <= 32'hfa6484bb;
			S3[126] <= 32'h8d6612ae; S3[127] <= 32'hbf3c6f47; S3[128] <= 32'hd29be463; 
			S3[129] <= 32'h542f5d9e; S3[130] <= 32'haec2771b; S3[131] <= 32'hf64e6370;
			S3[132] <= 32'h740e0d8d; S3[133] <= 32'he75b1357; S3[134] <= 32'hf8721671; 
			S3[135] <= 32'haf537d5d; S3[136] <= 32'h4040cb08; S3[137] <= 32'h4eb4e2cc;
			S3[138] <= 32'h34d2466a; S3[139] <= 32'h0115af84; S3[140] <= 32'he1b00428; 
			S3[141] <= 32'h95983a1d; S3[142] <= 32'h06b89fb4; S3[143] <= 32'hce6ea048;
			S3[144] <= 32'h6f3f3b82; S3[145] <= 32'h3520ab82; S3[146] <= 32'h011a1d4b; 
			S3[147] <= 32'h277227f8; S3[148] <= 32'h611560b1; S3[149] <= 32'he7933fdc;
			S3[150] <= 32'hbb3a792b; S3[151] <= 32'h344525bd; S3[152] <= 32'ha08839e1; 
			S3[153] <= 32'h51ce794b; S3[154] <= 32'h2f32c9b7; S3[155] <= 32'ha01fbac9;
			S3[156] <= 32'he01cc87e; S3[157] <= 32'hbcc7d1f6; S3[158] <= 32'hcf0111c3; 
			S3[159] <= 32'ha1e8aac7; S3[160] <= 32'h1a908749; S3[161] <= 32'hd44fbd9a;
			S3[162] <= 32'hd0dadecb; S3[163] <= 32'hd50ada38; S3[164] <= 32'h0339c32a; 
			S3[165] <= 32'hc6913667; S3[166] <= 32'h8df9317c; S3[167] <= 32'he0b12b4f;
			S3[168] <= 32'hf79e59b7; S3[169] <= 32'h43f5bb3a; S3[170] <= 32'hf2d519ff; 
			S3[171] <= 32'h27d9459c; S3[172] <= 32'hbf97222c; S3[173] <= 32'h15e6fc2a;
			S3[174] <= 32'h0f91fc71; S3[175] <= 32'h9b941525; S3[176] <= 32'hfae59361; 
			S3[177] <= 32'hceb69ceb; S3[178] <= 32'hc2a86459; S3[179] <= 32'h12baa8d1;
			S3[180] <= 32'hb6c1075e; S3[181] <= 32'he3056a0c; S3[182] <= 32'h10d25065; 
			S3[183] <= 32'hcb03a442; S3[184] <= 32'he0ec6e0e; S3[185] <= 32'h1698db3b;
			S3[186] <= 32'h4c98a0be; S3[187] <= 32'h3278e964; S3[188] <= 32'h9f1f9532; 
			S3[189] <= 32'he0d392df; S3[190] <= 32'hd3a0342b; S3[191] <= 32'h8971f21e;
			S3[192] <= 32'h1b0a7441; S3[193] <= 32'h4ba3348c; S3[194] <= 32'hc5be7120; 
			S3[195] <= 32'hc37632d8; S3[196] <= 32'hdf359f8d; S3[197] <= 32'h9b992f2e;
			S3[198] <= 32'he60b6f47; S3[199] <= 32'h0fe3f11d; S3[200] <= 32'he54cda54; 
			S3[201] <= 32'h1edad891; S3[202] <= 32'hce6279cf; S3[203] <= 32'hcd3e7e6f;
			S3[204] <= 32'h1618b166; S3[205] <= 32'hfd2c1d05; S3[206] <= 32'h848fd2c5; 
			S3[207] <= 32'hf6fb2299; S3[208] <= 32'hf523f357; S3[209] <= 32'ha6327623;
			S3[210] <= 32'h93a83531; S3[211] <= 32'h56cccd02; S3[212] <= 32'hacf08162; 
			S3[213] <= 32'h5a75ebb5; S3[214] <= 32'h6e163697; S3[215] <= 32'h88d273cc;
			S3[216] <= 32'hde966292; S3[217] <= 32'h81b949d0; S3[218] <= 32'h4c50901b; 
			S3[219] <= 32'h71c65614; S3[220] <= 32'he6c6c7bd; S3[221] <= 32'h327a140a;
			S3[222] <= 32'h45e1d006; S3[223] <= 32'hc3f27b9a; S3[224] <= 32'hc9aa53fd; 
			S3[225] <= 32'h62a80f00; S3[226] <= 32'hbb25bfe2; S3[227] <= 32'h35bdd2f6;
			S3[228] <= 32'h71126905; S3[229] <= 32'hb2040222; S3[230] <= 32'hb6cbcf7c; 
			S3[231] <= 32'hcd769c2b; S3[232] <= 32'h53113ec0; S3[233] <= 32'h1640e3d3;
			S3[234] <= 32'h38abbd60; S3[235] <= 32'h2547adf0; S3[236] <= 32'hba38209c; 
			S3[237] <= 32'hf746ce76; S3[238] <= 32'h77afa1c5; S3[239] <= 32'h20756060;
			S3[240] <= 32'h85cbfe4e; S3[241] <= 32'h8ae88dd8; S3[242] <= 32'h7aaaf9b0; 
			S3[243] <= 32'h4cf9aa7e; S3[244] <= 32'h1948c25c; S3[245] <= 32'h02fb8a8c;
			S3[246] <= 32'h01c36ae4; S3[247] <= 32'hd6ebe1f9; S3[248] <= 32'h90d4f869; 
			S3[249] <= 32'ha65cdea0; S3[250] <= 32'h3f09252d; S3[251] <= 32'hc208e69f;
			S3[252] <= 32'hb74e6132; S3[253] <= 32'hce77e25b; S3[254] <= 32'h578fdfe3; 
			S3[255] <= 32'h3ac372e6;

			initDone <= 1'b1;
			
		end
		
		else if(initDone)
		begin
			expandKey(Salt, Key);
			for (q = 0; q < cost - 1; q = q+1)
			begin
				for (y = 0; y < cost - 1; y = y+1)
				begin
					expandKey(128'd0, Key);
					expandKey(128'd0, {Salt, Salt, Salt, Salt, Salt[127:64]});
				end
			end
			expandDone = 0;
			
		end
		
		else if(expandDone)
		begin
			for (ecb = 0; ecb < 64; ecb = ecb + 1)
			begin
				cyph[191:128] = Encrypt(cyph[191:128]);
				cyph[127:64] = Encrypt(cyph[127:64]);
				cyph[63:0] = Encrypt(cyph[63:0]);
			end
			cryptmw <= {cost, Salt, cyph};
		end
		
	end
	assign cryptm = cryptmw;
endmodule
